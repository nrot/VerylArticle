module hello_Hello ();
    initial begin
        $display("hello world");
    end
endmodule
