module hello_ModuleA #(
    parameter int unsigned A = 10 ,
    parameter string       B = "" ,
    parameter int signed   C = -10,
    parameter int unsigned D = 0  
) (
    input logic clk
);

endmodule
